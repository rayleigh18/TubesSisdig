LIBRARY  IEEE; 
USE  IEEE.STD_LOGIC_1164.ALL; 
USE  IEEE.STD_LOGIC_ARITH.ALL; 
USE  IEEE.STD_LOGIC_UNSIGNED.ALL;
entity p1Win is
	port(
		x, y, rgb : in integer;
		outRGB    : out integer;
	);
end p1Win;

architecture structural of p1Win is

begin

image1(0,0,0) <= 99;
image1(0,0,1) <= 30;
image1(0,0,2) <= 233;
image1(0,1,0) <= 99;
image1(0,1,1) <= 30;
image1(0,1,2) <= 233;
image1(0,2,0) <= 99;
image1(0,2,1) <= 30;
image1(0,2,2) <= 233;
image1(0,3,0) <= 0;
image1(0,3,1) <= 0;
image1(0,3,2) <= 0;
image1(0,4,0) <= 0;
image1(0,4,1) <= 0;
image1(0,4,2) <= 0;
image1(1,0,0) <= 99;
image1(1,0,1) <= 30;
image1(1,0,2) <= 233;
image1(1,1,0) <= 0;
image1(1,1,1) <= 0;
image1(1,1,2) <= 0;
image1(1,2,0) <= 0;
image1(1,2,1) <= 0;
image1(1,2,2) <= 0;
image1(1,3,0) <= 99;
image1(1,3,1) <= 30;
image1(1,3,2) <= 233;
image1(1,4,0) <= 0;
image1(1,4,1) <= 0;
image1(1,4,2) <= 0;
image1(2,0,0) <= 99;
image1(2,0,1) <= 30;
image1(2,0,2) <= 233;
image1(2,1,0) <= 99;
image1(2,1,1) <= 30;
image1(2,1,2) <= 233;
image1(2,2,0) <= 99;
image1(2,2,1) <= 30;
image1(2,2,2) <= 233;
image1(2,3,0) <= 0;
image1(2,3,1) <= 0;
image1(2,3,2) <= 0;
image1(2,4,0) <= 0;
image1(2,4,1) <= 0;
image1(2,4,2) <= 0;
image1(3,0,0) <= 99;
image1(3,0,1) <= 30;
image1(3,0,2) <= 233;
image1(3,1,0) <= 0;
image1(3,1,1) <= 0;
image1(3,1,2) <= 0;
image1(3,2,0) <= 0;
image1(3,2,1) <= 0;
image1(3,2,2) <= 0;
image1(3,3,0) <= 0;
image1(3,3,1) <= 0;
image1(3,3,2) <= 0;
image1(3,4,0) <= 0;
image1(3,4,1) <= 0;
image1(3,4,2) <= 0;
image1(4,0,0) <= 99;
image1(4,0,1) <= 30;
image1(4,0,2) <= 233;
image1(4,1,0) <= 0;
image1(4,1,1) <= 0;
image1(4,1,2) <= 0;
image1(4,2,0) <= 0;
image1(4,2,1) <= 0;
image1(4,2,2) <= 0;
image1(4,3,0) <= 0;
image1(4,3,1) <= 0;
image1(4,3,2) <= 0;
image1(4,4,0) <= 0;
image1(4,4,1) <= 0;
image1(4,4,2) <= 0;
image1(5,0,0) <= 0;
image1(5,0,1) <= 0;
image1(5,0,2) <= 0;
image1(5,1,0) <= 0;
image1(5,1,1) <= 0;
image1(5,1,2) <= 0;
image1(5,2,0) <= 0;
image1(5,2,1) <= 0;
image1(5,2,2) <= 0;
image1(5,3,0) <= 0;
image1(5,3,1) <= 0;
image1(5,3,2) <= 0;
image1(5,4,0) <= 0;
image1(5,4,1) <= 0;
image1(5,4,2) <= 0;
image1(6,0,0) <= 0;
image1(6,0,1) <= 0;
image1(6,0,2) <= 0;
image1(6,1,0) <= 0;
image1(6,1,1) <= 0;
image1(6,1,2) <= 0;
image1(6,2,0) <= 0;
image1(6,2,1) <= 0;
image1(6,2,2) <= 0;
image1(6,3,0) <= 0;
image1(6,3,1) <= 0;
image1(6,3,2) <= 0;
image1(6,4,0) <= 0;
image1(6,4,1) <= 0;
image1(6,4,2) <= 0;
image1(7,0,0) <= 0;
image1(7,0,1) <= 0;
image1(7,0,2) <= 0;
image1(7,1,0) <= 0;
image1(7,1,1) <= 0;
image1(7,1,2) <= 0;
image1(7,2,0) <= 0;
image1(7,2,1) <= 0;
image1(7,2,2) <= 0;
image1(7,3,0) <= 0;
image1(7,3,1) <= 0;
image1(7,3,2) <= 0;
image1(7,4,0) <= 0;
image1(7,4,1) <= 0;
image1(7,4,2) <= 0;
image1(8,0,0) <= 0;
image1(8,0,1) <= 0;
image1(8,0,2) <= 0;
image1(8,1,0) <= 0;
image1(8,1,1) <= 0;
image1(8,1,2) <= 0;
image1(8,2,0) <= 0;
image1(8,2,1) <= 0;
image1(8,2,2) <= 0;
image1(8,3,0) <= 0;
image1(8,3,1) <= 0;
image1(8,3,2) <= 0;
image1(8,4,0) <= 0;
image1(8,4,1) <= 0;
image1(8,4,2) <= 0;
image1(9,0,0) <= 0;
image1(9,0,1) <= 0;
image1(9,0,2) <= 0;
image1(9,1,0) <= 0;
image1(9,1,1) <= 0;
image1(9,1,2) <= 0;
image1(9,2,0) <= 0;
image1(9,2,1) <= 0;
image1(9,2,2) <= 0;
image1(9,3,0) <= 0;
image1(9,3,1) <= 0;
image1(9,3,2) <= 0;
image1(9,4,0) <= 0;
image1(9,4,1) <= 0;
image1(9,4,2) <= 0;
image1(10,0,0) <= 0;
image1(10,0,1) <= 0;
image1(10,0,2) <= 0;
image1(10,1,0) <= 0;
image1(10,1,1) <= 0;
image1(10,1,2) <= 0;
image1(10,2,0) <= 0;
image1(10,2,1) <= 0;
image1(10,2,2) <= 0;
image1(10,3,0) <= 0;
image1(10,3,1) <= 0;
image1(10,3,2) <= 0;
image1(10,4,0) <= 0;
image1(10,4,1) <= 0;
image1(10,4,2) <= 0;
image1(11,0,0) <= 0;
image1(11,0,1) <= 0;
image1(11,0,2) <= 0;
image1(11,1,0) <= 0;
image1(11,1,1) <= 0;
image1(11,1,2) <= 0;
image1(11,2,0) <= 0;
image1(11,2,1) <= 0;
image1(11,2,2) <= 0;
image1(11,3,0) <= 0;
image1(11,3,1) <= 0;
image1(11,3,2) <= 0;
image1(11,4,0) <= 0;
image1(11,4,1) <= 0;
image1(11,4,2) <= 0;
image1(12,0,0) <= 0;
image1(12,0,1) <= 0;
image1(12,0,2) <= 0;
image1(12,1,0) <= 0;
image1(12,1,1) <= 0;
image1(12,1,2) <= 0;
image1(12,2,0) <= 0;
image1(12,2,1) <= 0;
image1(12,2,2) <= 0;
image1(12,3,0) <= 0;
image1(12,3,1) <= 0;
image1(12,3,2) <= 0;
image1(12,4,0) <= 0;
image1(12,4,1) <= 0;
image1(12,4,2) <= 0;
image1(13,0,0) <= 0;
image1(13,0,1) <= 0;
image1(13,0,2) <= 0;
image1(13,1,0) <= 0;
image1(13,1,1) <= 0;
image1(13,1,2) <= 0;
image1(13,2,0) <= 0;
image1(13,2,1) <= 0;
image1(13,2,2) <= 0;
image1(13,3,0) <= 0;
image1(13,3,1) <= 0;
image1(13,3,2) <= 0;
image1(13,4,0) <= 0;
image1(13,4,1) <= 0;
image1(13,4,2) <= 0;
image1(14,0,0) <= 0;
image1(14,0,1) <= 0;
image1(14,0,2) <= 0;
image1(14,1,0) <= 0;
image1(14,1,1) <= 0;
image1(14,1,2) <= 0;
image1(14,2,0) <= 0;
image1(14,2,1) <= 0;
image1(14,2,2) <= 0;
image1(14,3,0) <= 0;
image1(14,3,1) <= 0;
image1(14,3,2) <= 0;
image1(14,4,0) <= 0;
image1(14,4,1) <= 0;
image1(14,4,2) <= 0;
image1(15,0,0) <= 0;
image1(15,0,1) <= 0;
image1(15,0,2) <= 0;
image1(15,1,0) <= 0;
image1(15,1,1) <= 0;
image1(15,1,2) <= 0;
image1(15,2,0) <= 0;
image1(15,2,1) <= 0;
image1(15,2,2) <= 0;
image1(15,3,0) <= 0;
image1(15,3,1) <= 0;
image1(15,3,2) <= 0;
image1(15,4,0) <= 0;
image1(15,4,1) <= 0;
image1(15,4,2) <= 0;
image1(16,0,0) <= 0;
image1(16,0,1) <= 0;
image1(16,0,2) <= 0;
image1(16,1,0) <= 0;
image1(16,1,1) <= 0;
image1(16,1,2) <= 0;
image1(16,2,0) <= 0;
image1(16,2,1) <= 0;
image1(16,2,2) <= 0;
image1(16,3,0) <= 0;
image1(16,3,1) <= 0;
image1(16,3,2) <= 0;
image1(16,4,0) <= 0;
image1(16,4,1) <= 0;
image1(16,4,2) <= 0;
image1(17,0,0) <= 0;
image1(17,0,1) <= 0;
image1(17,0,2) <= 0;
image1(17,1,0) <= 0;
image1(17,1,1) <= 0;
image1(17,1,2) <= 0;
image1(17,2,0) <= 0;
image1(17,2,1) <= 0;
image1(17,2,2) <= 0;
image1(17,3,0) <= 0;
image1(17,3,1) <= 0;
image1(17,3,2) <= 0;
image1(17,4,0) <= 0;
image1(17,4,1) <= 0;
image1(17,4,2) <= 0;
image1(18,0,0) <= 0;
image1(18,0,1) <= 0;
image1(18,0,2) <= 0;
image1(18,1,0) <= 0;
image1(18,1,1) <= 0;
image1(18,1,2) <= 0;
image1(18,2,0) <= 0;
image1(18,2,1) <= 0;
image1(18,2,2) <= 0;
image1(18,3,0) <= 0;
image1(18,3,1) <= 0;
image1(18,3,2) <= 0;
image1(18,4,0) <= 0;
image1(18,4,1) <= 0;
image1(18,4,2) <= 0;
image1(19,0,0) <= 0;
image1(19,0,1) <= 0;
image1(19,0,2) <= 0;
image1(19,1,0) <= 0;
image1(19,1,1) <= 0;
image1(19,1,2) <= 0;
image1(19,2,0) <= 0;
image1(19,2,1) <= 0;
image1(19,2,2) <= 0;
image1(19,3,0) <= 0;
image1(19,3,1) <= 0;
image1(19,3,2) <= 0;
image1(19,4,0) <= 0;
image1(19,4,1) <= 0;
image1(19,4,2) <= 0;
image1(20,0,0) <= 0;
image1(20,0,1) <= 0;
image1(20,0,2) <= 0;
image1(20,1,0) <= 0;
image1(20,1,1) <= 0;
image1(20,1,2) <= 0;
image1(20,2,0) <= 0;
image1(20,2,1) <= 0;
image1(20,2,2) <= 0;
image1(20,3,0) <= 0;
image1(20,3,1) <= 0;
image1(20,3,2) <= 0;
image1(20,4,0) <= 0;
image1(20,4,1) <= 0;
image1(20,4,2) <= 0;
image1(21,0,0) <= 0;
image1(21,0,1) <= 0;
image1(21,0,2) <= 0;
image1(21,1,0) <= 0;
image1(21,1,1) <= 0;
image1(21,1,2) <= 0;
image1(21,2,0) <= 0;
image1(21,2,1) <= 0;
image1(21,2,2) <= 0;
image1(21,3,0) <= 0;
image1(21,3,1) <= 0;
image1(21,3,2) <= 0;
image1(21,4,0) <= 0;
image1(21,4,1) <= 0;
image1(21,4,2) <= 0;
image1(22,0,0) <= 0;
image1(22,0,1) <= 0;
image1(22,0,2) <= 0;
image1(22,1,0) <= 0;
image1(22,1,1) <= 0;
image1(22,1,2) <= 0;
image1(22,2,0) <= 0;
image1(22,2,1) <= 0;
image1(22,2,2) <= 0;
image1(22,3,0) <= 0;
image1(22,3,1) <= 0;
image1(22,3,2) <= 0;
image1(22,4,0) <= 0;
image1(22,4,1) <= 0;
image1(22,4,2) <= 0;
image1(23,0,0) <= 0;
image1(23,0,1) <= 0;
image1(23,0,2) <= 0;
image1(23,1,0) <= 0;
image1(23,1,1) <= 0;
image1(23,1,2) <= 0;
image1(23,2,0) <= 0;
image1(23,2,1) <= 0;
image1(23,2,2) <= 0;
image1(23,3,0) <= 0;
image1(23,3,1) <= 0;
image1(23,3,2) <= 0;
image1(23,4,0) <= 0;
image1(23,4,1) <= 0;
image1(23,4,2) <= 0;
image1(24,0,0) <= 0;
image1(24,0,1) <= 0;
image1(24,0,2) <= 0;
image1(24,1,0) <= 0;
image1(24,1,1) <= 0;
image1(24,1,2) <= 0;
image1(24,2,0) <= 0;
image1(24,2,1) <= 0;
image1(24,2,2) <= 0;
image1(24,3,0) <= 0;
image1(24,3,1) <= 0;
image1(24,3,2) <= 0;
image1(24,4,0) <= 0;
image1(24,4,1) <= 0;
image1(24,4,2) <= 0;
